module and_gate_s(a,b,y);
input a,b;
output y;

and(y,a,b);
                
endmodule